`timescale 1ns/1ns

module write_memory;

endmodule